module main

fn test_input() {
	assert defrag('input_test.txt') == 1928
}
