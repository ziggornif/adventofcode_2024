module main

fn test_input() {
	assert antinodes('input_test.txt') == 14
}
